



module testFullAdder();

   reg [2:0] switches;

   wire 